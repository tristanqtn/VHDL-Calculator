-- LIBRAIRIES ----------------------------------------------------------------------------
LIBRARY IEEE;
USE work.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
------------------------------------------------------------------------------------------

------------------------------------------------------------------------------------------
-- AFFICHAGE -----------------------------------------------------------------------------
------------------------------------------------------------------------------------------
ENTITY affichage IS

	PORT (
		resultat : IN std_logic_vector (7 DOWNTO 0); -- choix du type d'opération à effectuer (2 bits)
		signe : IN std_logic;
 
		seg1, seg2, seg3, seg4 : OUT std_logic_vector(7 DOWNTO 0) -- chaque variable correspond à un afficheur 7seg (8 bits)
	);
 
END affichage;
------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------


------------------------------------------------------------------------------------------
--ARCHITECTURE DE L4AFFICHAGE ------------------------------------------------------------
------------------------------------------------------------------------------------------
ARCHITECTURE bhv OF affichage IS

	SIGNAL c : std_logic_vector(7 DOWNTO 0);

BEGIN
	PROCESS (resultat) -- dès qu'un changment d'etat est repéré sur resultat
	BEGIN
		c <= resultat; --stockage du resulatat unsigned dnas le signal temporaire c
 
		IF (c(7) = '1' AND signe = '1') THEN
			seg4 <= "10111111";
		ELSE
			seg4 <= "11111111";
		END IF;
 
		IF (signe = '1') THEN
			IF (c(6 DOWNTO 0) = "0000000") THEN -- 0 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0000001") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0000010") THEN --2
				seg1 <= "10100100";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0000011") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0000100") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0000101") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0000110") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0000111") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0001000") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0001001") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0001010") THEN -- 0 10 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0001011") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0001100") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0001101") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0001110") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0001111") THEN -- 5 
				seg1 <= "10010010";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0010000") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0010001") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0010010") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0010011") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0010100") THEN -- 0 20 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0010101") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0010110") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0010111") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0011000") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0011001") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0011010") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0011011") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0011100") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0011101") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0011110") THEN -- 0 30 ------------------------------------------- 
				seg1 <= "11000000"; 
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0011111") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0100000") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0100001") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0100010") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0100011") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0100100") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0100101") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0100110") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0100111") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0101000") THEN -- 0 40 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0101001") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0101010") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0101011") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0101100") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0101101") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0101110") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0101111") THEN -- 7 
				seg1 <= "11111000";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0110000") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c(6 DOWNTO 0) = "0110001") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10011001";
				seg3 <= "11000000"; --50 -------------------------------------------
			END IF;
 
		ELSE
 
			IF (c = "00000000") THEN -- 0 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c = "00000001") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c = "00000010") THEN --2
				seg1 <= "10100100";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c = "00000011") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c = "00000100") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c = "00000101") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c = "00000110") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c = "00000111") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c = "00001000") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c = "00001001") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "11000000";
				seg3 <= "11000000";
			ELSIF (c = "00001010") THEN -- 0 10 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c = "00001011") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c = "00001100") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c = "00001101") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c = "00001110") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c = "00001111") THEN -- 5 
				seg1 <= "10010010";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c = "00010000") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c = "00010001") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c = "00010010") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c = "00010011") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "11111001";
				seg3 <= "11000000";
			ELSIF (c = "00010100") THEN -- 0 20 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c = "00010101") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c = "00010110") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c = "00010111") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c = "00011000") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c = "00011001") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c = "00011010") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c = "00011011") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c = "00011100") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c = "00011101") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10100100";
				seg3 <= "11000000";
			ELSIF (c = "00011110") THEN -- 0 30 ------------------------------------------- 
				seg1 <= "11000000"; 
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c = "00011111") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c = "00100000") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c = "00100001") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c = "00100010") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c = "00100011") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c = "00100100") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c = "00100101") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c = "00100110") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c = "00100111") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10110000";
				seg3 <= "11000000";
			ELSIF (c = "00101000") THEN -- 0 40 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c = "00101001") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c = "00101010") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c = "00101011") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c = "00101100") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c = "00101101") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c = "00101110") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c = "00101111") THEN -- 7 
				seg1 <= "11111000";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c = "00110000") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10011001";
				seg3 <= "11000000";
			ELSIF (c = "00110001") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10011001";
				seg3 <= "11000000"; --50 -------------------------------------------
			ELSIF (c = "00110010") THEN -- 0
				seg1 <= "11000000"; 
				seg2 <= "10010010";
				seg3 <= "11000000";
			ELSIF (c = "00110011") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10010010";
				seg3 <= "11000000";
			ELSIF (c = "00110100") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10010010";
				seg3 <= "11000000";
			ELSIF (c = "00110101") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10010010";
				seg3 <= "11000000";
			ELSIF (c = "00110110") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10010010";
				seg3 <= "11000000";
			ELSIF (c = "00110111") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10010010";
				seg3 <= "11000000";
			ELSIF (c = "00111000") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10010010";
				seg3 <= "11000000";
			ELSIF (c = "00111001") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10010010";
				seg3 <= "11000000";
			ELSIF (c = "00111010") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10010010";
				seg3 <= "11000000";
			ELSIF (c = "00111011") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10010010";
				seg3 <= "11000000";
			ELSIF (c = "00111100") THEN -- 0 60 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10000010";
				seg3 <= "11000000";
			ELSIF (c = "00111101") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10000010";
				seg3 <= "11000000";
			ELSIF (c = "00111110") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10000010";
				seg3 <= "11000000";
			ELSIF (c = "00111111") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10000010";
				seg3 <= "11000000";
			ELSIF (c = "01000000") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10000010";
				seg3 <= "11000000";
			ELSIF (c = "01000001") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10000010";
				seg3 <= "11000000";
			ELSIF (c = "01000010") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10000010";
				seg3 <= "11000000";
			ELSIF (c = "01000011") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10000010";
				seg3 <= "11000000";
			ELSIF (c = "01000100") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10000010";
				seg3 <= "11000000";
			ELSIF (c = "01000101") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10000010";
				seg3 <= "11000000";
			ELSIF (c = "01000110") THEN -- 0 70 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "11111000";
				seg3 <= "11000000";
			ELSIF (c = "01000111") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "11111000";
				seg3 <= "11000000";
			ELSIF (c = "01001000") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "11111000";
				seg3 <= "11000000";
			ELSIF (c = "01001001") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "11111000";
				seg3 <= "11000000";
			ELSIF (c = "01001010") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "11111000";
				seg3 <= "11000000";
			ELSIF (c = "01001011") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "11111000";
				seg3 <= "11000000";
			ELSIF (c = "01001100") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "11111000";
				seg3 <= "11000000";
			ELSIF (c = "01001101") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "11111000";
				seg3 <= "11000000";
			ELSIF (c = "01001110") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "11111000";
				seg3 <= "11000000";
			ELSIF (c = "01001111") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "11111000";
				seg3 <= "11000000";
			ELSIF (c = "01010000") THEN -- 0 80 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10000000";
				seg3 <= "11000000";
			ELSIF (c = "01010001") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10000000";
				seg3 <= "11000000";
			ELSIF (c = "01010010") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10000000";
				seg3 <= "11000000";
			ELSIF (c = "01010011") THEN -- 3 
				seg1 <= "10110000";
				seg2 <= "10000000";
				seg3 <= "11000000";
			ELSIF (c = "01010100") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10000000";
				seg3 <= "11000000";
			ELSIF (c = "01010101") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10000000";
				seg3 <= "11000000";
			ELSIF (c = "01010110") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10000000";
				seg3 <= "11000000";
			ELSIF (c = "01010111") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10000000";
				seg3 <= "11000000";
			ELSIF (c = "01011000") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10000000";
				seg3 <= "11000000";
			ELSIF (c = "01011001") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10000000";
				seg3 <= "11000000";
			ELSIF (c = "01011010") THEN -- 0 90 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10010000";
				seg3 <= "11000000";
			ELSIF (c = "01011011") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10010000";
				seg3 <= "11000000";
			ELSIF (c = "01011100") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10010000";
				seg3 <= "11000000";
			ELSIF (c = "01011101") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10010000";
				seg3 <= "11000000";
			ELSIF (c = "01011110") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10010000";
				seg3 <= "11000000";
			ELSIF (c = "01011111") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10010000";
				seg3 <= "11000000";
			ELSIF (c = "01100000") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10010000";
				seg3 <= "11000000";
			ELSIF (c = "01100001") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10010000";
				seg3 <= "11000000";
			ELSIF (c = "01100010") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10010000";
				seg3 <= "11000000";
			ELSIF (c = "01100011") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10010000";
				seg3 <= "11000000"; 
			ELSIF (c = "01100100") THEN -- 0 100 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "11000000";
				seg3 <= "11111001";
			ELSIF (c = "01100101") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "11000000";
				seg3 <= "11111001";
			ELSIF (c = "01100110") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "11000000";
				seg3 <= "11111001";
			ELSIF (c = "01100111") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "11000000";
				seg3 <= "11111001";
			ELSIF (c = "01101000") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "11000000";
				seg3 <= "11111001";
			ELSIF (c = "01101001") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "11000000";
				seg3 <= "11111001";
			ELSIF (c = "01101010") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "11000000";
				seg3 <= "11111001";
			ELSIF (c = "01101011") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "11000000";
				seg3 <= "11111001";
			ELSIF (c = "01101100") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "11000000";
				seg3 <= "11111001";
			ELSIF (c = "01101101") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "11000000";
				seg3 <= "11111001";
			ELSIF (c = "01101110") THEN -- 0 110 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "11111001";
				seg3 <= "11111001";
			ELSIF (c = "01101111") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "11111001";
				seg3 <= "11111001";
			ELSIF (c = "01110000") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "11111001";
				seg3 <= "11111001";
			ELSIF (c = "01110001") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "11111001";
				seg3 <= "11111001";
			ELSIF (c = "01110010") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "11111001";
				seg3 <= "11111001";
			ELSIF (c = "01110011") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10010010";
				seg3 <= "11111001";
			ELSIF (c = "01110100") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "11111001";
				seg3 <= "11111001";
			ELSIF (c = "01110101") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "11111001";
				seg3 <= "11111001";
			ELSIF (c = "01110110") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "11111001";
				seg3 <= "11111001";
			ELSIF (c = "01110111") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "11111001";
				seg3 <= "11111001";
			ELSIF (c = "01111000") THEN -- 0 120 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10100100";
				seg3 <= "11111001";
			ELSIF (c = "01111001") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10100100";
				seg3 <= "11111001";
			ELSIF (c = "01111010") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10100100";
				seg3 <= "11111001";
			ELSIF (c = "01111011") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10100100";
				seg3 <= "11111001";
			ELSIF (c = "01111100") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10100100";
				seg3 <= "11111001";
			ELSIF (c = "01111101") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10100100";
				seg3 <= "11111001";
			ELSIF (c = "01111110") THEN -- 6 
				seg1 <= "10000010";
				seg2 <= "10100100";
				seg3 <= "11111001";
			ELSIF (c = "01111111") THEN -- 7 
				seg1 <= "11111000";
				seg2 <= "10100100";
				seg3 <= "11111001";
			ELSIF (c = "10000000") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10100100";
				seg3 <= "11111001";
			ELSIF (c = "10000001") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10100100";
				seg3 <= "11111001";
			ELSIF (c = "10000010") THEN -- 0 130 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10110000";
				seg3 <= "11111001";
			ELSIF (c = "10000011") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10110000";
				seg3 <= "11111001";
			ELSIF (c = "10000100") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10110000";
				seg3 <= "11111001";
			ELSIF (c = "10000101") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10110000";
				seg3 <= "11111001";
			ELSIF (c = "10000110") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10110000";
				seg3 <= "11111001";
			ELSIF (c = "10000111") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10110000";
				seg3 <= "11111001";
			ELSIF (c = "10001000") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10110000";
				seg3 <= "11111001";
			ELSIF (c = "10001001") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10110000";
				seg3 <= "11111001";
			ELSIF (c = "10001010") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10110000";
				seg3 <= "11111001";
			ELSIF (c = "10001011") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10110000";
				seg3 <= "11111001";
			ELSIF (c = "10001100") THEN -- 0 140 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10011001";
				seg3 <= "11111001";
			ELSIF (c = "10001101") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10011001";
				seg3 <= "11111001";
			ELSIF (c = "10001110") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10011001";
				seg3 <= "11111001";
			ELSIF (c = "10001111") THEN -- 3 
				seg1 <= "10110000";
				seg2 <= "10011001";
				seg3 <= "11111001";
			ELSIF (c = "10010000") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10011001";
				seg3 <= "11111001";
			ELSIF (c = "10010001") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10011001";
				seg3 <= "11111001";
			ELSIF (c = "10010010") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10011001";
				seg3 <= "11111001";
			ELSIF (c = "10010011") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10011001";
				seg3 <= "11111001";
			ELSIF (c = "10010100") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10011001";
				seg3 <= "11111001";
			ELSIF (c = "10010101") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10011001";
				seg3 <= "11111001"; 
			ELSIF (c = "10010110") THEN -- 0 150 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10010010";
				seg3 <= "11111001";
			ELSIF (c = "10010111") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10010010";
				seg3 <= "11111001";
			ELSIF (c = "10011000") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10010010";
				seg3 <= "11111001";
			ELSIF (c = "10011001") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10010010";
				seg3 <= "11111001";
			ELSIF (c = "10011010") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10010010";
				seg3 <= "11111001";
			ELSIF (c = "10011011") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10010010";
				seg3 <= "11111001";
			ELSIF (c = "10011100") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10010010";
				seg3 <= "11111001";
			ELSIF (c = "10011101") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10010010";
				seg3 <= "11111001";
			ELSIF (c = "10011110") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10010010";
				seg3 <= "11111001";
			ELSIF (c = "10011111") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10010010";
				seg3 <= "11111001";
			ELSIF (c = "10100000") THEN -- 0 160 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10000010";
				seg3 <= "11111001";
			ELSIF (c = "10100001") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10000010";
				seg3 <= "11111001";
			ELSIF (c = "10100010") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10000010";
				seg3 <= "11111001";
			ELSIF (c = "10100011") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10000010";
				seg3 <= "11111001";
			ELSIF (c = "10100100") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10000010";
				seg3 <= "11111001";
			ELSIF (c = "10100101") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10000010";
				seg3 <= "11111001";
			ELSIF (c = "10100110") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10000010";
				seg3 <= "11111001";
			ELSIF (c = "10100111") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10000010";
				seg3 <= "11111001";
			ELSIF (c = "10101000") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10000010";
				seg3 <= "11111001";
			ELSIF (c = "10101001") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10000010";
				seg3 <= "11111001";
			ELSIF (c = "10101010") THEN -- 0 170 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "11111000";
				seg3 <= "11111001";
			ELSIF (c = "10101011") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "11111000";
				seg3 <= "11111001";
			ELSIF (c = "10101100") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "11111000";
				seg3 <= "11111001";
			ELSIF (c = "10101101") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "11111000";
				seg3 <= "11111001";
			ELSIF (c = "10101110") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "11111000";
				seg3 <= "11111001";
			ELSIF (c = "10101111") THEN -- 5 
				seg1 <= "10010010";
				seg2 <= "11111000";
				seg3 <= "11111001";
			ELSIF (c = "10110000") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "11111000";
				seg3 <= "11111001";
			ELSIF (c = "10110001") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "11111000";
				seg3 <= "11111001";
			ELSIF (c = "10110010") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "11111000";
				seg3 <= "11111001";
			ELSIF (c = "10110011") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "11111000";
				seg3 <= "11111001";
			ELSIF (c = "10110100") THEN -- 0 180 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10000000";
				seg3 <= "11111001";
			ELSIF (c = "10110101") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10000000";
				seg3 <= "11111001";
			ELSIF (c = "10110110") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10000000";
				seg3 <= "11111001";
			ELSIF (c = "10110111") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10000000";
				seg3 <= "11111001";
			ELSIF (c = "10111000") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10000000";
				seg3 <= "11111001";
			ELSIF (c = "10111001") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10000000";
				seg3 <= "11111001";
			ELSIF (c = "10111010") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10000000";
				seg3 <= "11111001";
			ELSIF (c = "10111011") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10000000";
				seg3 <= "11111001";
			ELSIF (c = "10111100") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10000000";
				seg3 <= "11111001";
			ELSIF (c = "10111101") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10000000";
				seg3 <= "11111001";
			ELSIF (c = "10111110") THEN -- 0 190 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10010000";
				seg3 <= "11111001";
			ELSIF (c = "10111111") THEN -- 1 
				seg1 <= "11111001";
				seg2 <= "10010000";
				seg3 <= "11111001";
			ELSIF (c = "11000000") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10010000";
				seg3 <= "11111001";
			ELSIF (c = "11000001") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10010000";
				seg3 <= "11111001";
			ELSIF (c = "11000010") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10010000";
				seg3 <= "11111001";
			ELSIF (c = "11000011") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "10010000";
				seg3 <= "11111001";
			ELSIF (c = "11000100") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "10010000";
				seg3 <= "11111001";
			ELSIF (c = "11000101") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "10010000";
				seg3 <= "11111001";
			ELSIF (c = "11000110") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "10010000";
				seg3 <= "11111001";
			ELSIF (c = "11000111") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "10010000";
				seg3 <= "11111001"; 
			ELSIF (c = "11001000") THEN -- 0 200 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "11000000";
				seg3 <= "10100100";
			ELSIF (c = "11001001") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "11000000";
				seg3 <= "10100100";
			ELSIF (c = "11001010") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "11000000";
				seg3 <= "10100100";
			ELSIF (c = "11001011") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "11000000";
				seg3 <= "10100100";
			ELSIF (c = "11001100") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "11000000";
				seg3 <= "10100100";
			ELSIF (c = "11001101") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "11000000";
				seg3 <= "10100100";
			ELSIF (c = "11001110") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "11000000";
				seg3 <= "10100100";
			ELSIF (c = "11001111") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "11000000";
				seg3 <= "10100100";
			ELSIF (c = "11010000") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "11000000";
				seg3 <= "10100100";
			ELSIF (c = "11010001") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "11000000";
				seg3 <= "10100100";
			ELSIF (c = "11010010") THEN -- 0 210 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "11111001";
				seg3 <= "10100100";
			ELSIF (c = "11010011") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "11111001";
				seg3 <= "10100100";
			ELSIF (c = "11010100") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "11111001";
				seg3 <= "10100100";
			ELSIF (c = "11010101") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "11111001";
				seg3 <= "10100100";
			ELSIF (c = "11010110") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "11111001";
				seg3 <= "10100100";
			ELSIF (c = "11010111") THEN -- 5
				seg1 <= "10010010";
				seg2 <= "11111001";
				seg3 <= "10100100";
			ELSIF (c = "11011000") THEN -- 6
				seg1 <= "10000010";
				seg2 <= "11111001";
				seg3 <= "10100100";
			ELSIF (c = "11011001") THEN -- 7
				seg1 <= "11111000";
				seg2 <= "11111001";
				seg3 <= "10100100";
			ELSIF (c = "11011010") THEN -- 8
				seg1 <= "10000000";
				seg2 <= "11111001";
				seg3 <= "10100100";
			ELSIF (c = "11011011") THEN -- 9
				seg1 <= "10010000";
				seg2 <= "11111001";
				seg3 <= "10100100"; 
			ELSIF (c = "11011100") THEN -- 0 220 -------------------------------------------
				seg1 <= "11000000"; 
				seg2 <= "10100100";
				seg3 <= "10100100";
			ELSIF (c = "11011101") THEN -- 1
				seg1 <= "11111001";
				seg2 <= "10100100";
				seg3 <= "10100100";
			ELSIF (c = "11011110") THEN -- 2
				seg1 <= "10100100";
				seg2 <= "10100100";
				seg3 <= "10100100";
			ELSIF (c = "11011111") THEN -- 3
				seg1 <= "10110000";
				seg2 <= "10100100";
				seg3 <= "10100100";
			ELSIF (c = "11100000") THEN -- 4
				seg1 <= "10011001";
				seg2 <= "10100100";
				seg3 <= "10100100"; 
			ELSIF (c = "11100001") THEN -- 225 -------------------------------------------
				seg1 <= "10010010";
				seg2 <= "10100100";
				seg3 <= "10100100";
			END IF;
		END IF; -- fin du if
	END PROCESS; --fin du process
END bhv;
------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------