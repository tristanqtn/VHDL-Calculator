-- LIBRAIRIES ----------------------------------------------------------------------------
library IEEE;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
------------------------------------------------------------------------------------------



------------------------------------------------------------------------------------------
-- OPERATION NON SIGNEE ------------------------------------------------------------------
------------------------------------------------------------------------------------------
entity un_operation is 

    port( 
			 choix_op: in std_logic_vector (1 downto 0); -- choix du type d'opération à effectuer (2 bits)
		    operande_1, operande_2 : in std_logic_vector(3 downto 0); -- les deux opérandes reçues (4 bits)
			 
			 led_off : out std_logic_vector(1 downto 0); -- variable permettant d'eteindre les leds en trop (2 bits)
			 full_result : out std_logic_vector (7 downto 0); -- sortie de l'opération (8 bits)
			 seg1, seg2, seg3 : OUT std_logic_vector(7 downto 0) -- chaque variable correspond à un afficheur 7seg (8 bits)
		  );
		  
end un_operation; 
------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------


------------------------------------------------------------------------------------------
-- STRUCTURE OPERATION NON SIGNEE --------------------------------------------------------
------------------------------------------------------------------------------------------
architecture behavioral of un_operation is 

    signal un_result, sum, div, mult, sub, c : unsigned (7 downto 0); -- signaux utilisés pour les calculs 

begin

	sum <= unsigned("0000" & operande_1) + unsigned("0000" & operande_2); -- somme de deux vecteurs binaires non singés sur 4 bits 
	div <= "00000000" when unsigned(operande_2) = "0000" else (unsigned("0000" & operande_1) / unsigned("0000" & operande_2)); -- division euclidienne de deux vecteurs binaires non singés sur 4 bits si l'operande 2 n'est pas égale à 0000
	mult <= unsigned(operande_1) * unsigned(operande_2); -- multiplication de deux vecteurs binaires non singés sur 4 bits
	sub <= unsigned("0000" & operande_1) - unsigned("0000" & operande_2) when (unsigned(operande_1) >= unsigned(operande_2)) else "00000000"; -- différence dans les entiers naturels de deux vecteurs binaires non singés sur 4 bits
	
	--eteindre les leds inutilisées
	led_off(1) <= '0';
	led_off(0) <= '0';
	
	--sélection du résultat selon le type d'opération choisie
	WITH choix_op SELECT 

			un_result <= 	sum  when "00",
								mult when "10",
								sub  when "01",
								div  when "11";
			
    
	--stockage du résultat dans la sortie de l'entitée
	full_result <= std_logic_vector(un_result (7 downto 0));
	
	
	process(un_result) -- dès qu'un changment d'etat est repéré sur un_result
	begin
	
		c <= un_result; --stockage du resulatat unsigned dnas le signal temporaire c 
		
		
		if(c = "00000000")then	-- 0 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "11000000";
			seg3 <= "11000000";
		elsif(c = "00000001")then	-- 1
			seg1 <= "11111001";
			seg2 <= "11000000";
			seg3 <= "11000000";
		elsif(c = "00000010")then	--2
			seg1 <= "10100100";
			seg2 <= "11000000";
			seg3 <= "11000000";
		elsif(c = "00000011")then	-- 3
			seg1 <= "10110000";
			seg2 <= "11000000";
			seg3 <= "11000000";
		elsif(c = "00000100")then	-- 4
			seg1 <= "10011001";
			seg2 <= "11000000";
			seg3 <= "11000000";
		elsif(c = "00000101")then	-- 5
			seg1 <= "10010010";
			seg2 <= "11000000";
			seg3 <= "11000000";
		elsif(c = "00000110")then	-- 6
			seg1 <= "10000010";
			seg2 <= "11000000";
			seg3 <= "11000000";
		elsif(c = "00000111")then	-- 7
			seg1 <= "11111000";
			seg2 <= "11000000";
			seg3 <= "11000000";
		elsif(c = "00001000")then	-- 8
			seg1 <= "10000000";
			seg2 <= "11000000";
			seg3 <= "11000000";
		elsif(c = "00001001")then	-- 9
			seg1 <= "10010000";
			seg2 <= "11000000";
			seg3 <= "11000000";
		elsif(c = "00001010")then	-- 0	 10 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "11111001";
			seg3 <= "11000000";
		elsif(c = "00001011")then	-- 1
			seg1 <= "11111001";
			seg2 <= "11111001";
			seg3 <= "11000000";
		elsif(c = "00001100")then	-- 2
			seg1 <= "10100100";
			seg2 <= "11111001";
			seg3 <= "11000000";
		elsif(c = "00001101")then	-- 3
			seg1 <= "10110000";
			seg2 <= "11111001";
			seg3 <= "11000000";
		elsif(c = "00001110")then	-- 4
			seg1 <= "10011001";
			seg2 <= "11111001";
			seg3 <= "11000000";
		elsif(c = "00001111")then	-- 5	
			seg1 <= "10010010";
			seg2 <= "11111001";
			seg3 <= "11000000";
		elsif(c = "00010000")then	-- 6
			seg1 <= "10000010";
			seg2 <= "11111001";
			seg3 <= "11000000";
		elsif(c = "00010001")then	-- 7
			seg1 <= "11111000";
			seg2 <= "11111001";
			seg3 <= "11000000";
		elsif(c = "00010010")then	-- 8
			seg1 <= "10000000";
			seg2 <= "11111001";
			seg3 <= "11000000";
		elsif(c = "00010011")then	-- 9
			seg1 <= "10010000";
			seg2 <= "11111001";
			seg3 <= "11000000";
		elsif(c = "00010100")then	-- 0	20	-------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "10100100";
			seg3 <= "11000000";
		elsif(c = "00010101")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10100100";
			seg3 <= "11000000";
		elsif(c = "00010110")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10100100";
			seg3 <= "11000000";
		elsif(c = "00010111")then	-- 3
			seg1 <= "10110000";
			seg2 <= "10100100";
			seg3 <= "11000000";
		elsif(c = "00011000")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10100100";
			seg3 <= "11000000";
		elsif(c = "00011001")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10100100";
			seg3 <= "11000000";
		elsif(c = "00011010")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10100100";
			seg3 <= "11000000";
		elsif(c = "00011011")then	-- 7
			seg1 <= "11111000";
			seg2 <= "10100100";
			seg3 <= "11000000";
		elsif(c = "00011100")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10100100";
			seg3 <= "11000000";
		elsif(c = "00011101")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10100100";
			seg3 <= "11000000";
		elsif(c = "00011110")then	-- 0	30	-------------------------------------------	
			seg1 <= "11000000";	
			seg2 <= "10110000";
			seg3 <= "11000000";
		elsif(c = "00011111")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10110000";
			seg3 <= "11000000";
		elsif(c = "00100000")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10110000";
			seg3 <= "11000000";
		elsif(c = "00100001")then	-- 3
			seg1 <= "10110000";
			seg2 <= "10110000";
			seg3 <= "11000000";
		elsif(c = "00100010")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10110000";
			seg3 <= "11000000";
		elsif(c = "00100011")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10110000";
			seg3 <= "11000000";
		elsif(c = "00100100")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10110000";
			seg3 <= "11000000";
		elsif(c = "00100101")then	-- 7
			seg1 <= "11111000";
			seg2 <= "10110000";
			seg3 <= "11000000";
		elsif(c = "00100110")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10110000";
			seg3 <= "11000000";
		elsif(c = "00100111")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10110000";
			seg3 <= "11000000";
		elsif(c = "00101000")then	-- 0	40	-------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "10011001";
			seg3 <= "11000000";
		elsif(c = "00101001")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10011001";
			seg3 <= "11000000";
		elsif(c = "00101010")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10011001";
			seg3 <= "11000000";
		elsif(c = "00101011")then	-- 3
			seg1 <= "10110000";
			seg2 <= "10011001";
			seg3 <= "11000000";
		elsif(c = "00101100")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10011001";
			seg3 <= "11000000";
		elsif(c = "00101101")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10011001";
			seg3 <= "11000000";
		elsif(c = "00101110")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10011001";
			seg3 <= "11000000";
		elsif(c = "00101111")then	-- 7	
			seg1 <= "11111000";
			seg2 <= "10011001";
			seg3 <= "11000000";
		elsif(c = "00110000")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10011001";
			seg3 <= "11000000";
		elsif(c = "00110001")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10011001";
			seg3 <= "11000000";				--50 ------------------------------------------- 
		elsif(c = "00110010")then	-- 0
			seg1 <= "11000000";	
			seg2 <= "10010010";
			seg3 <= "11000000";
		elsif(c = "00110011")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10010010";
			seg3 <= "11000000";
		elsif(c = "00110100")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10010010";
			seg3 <= "11000000";
		elsif(c = "00110101")then	-- 3
			seg1 <= "10110000";
			seg2 <= "10010010";
			seg3 <= "11000000";
		elsif(c = "00110110")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10010010";
			seg3 <= "11000000";
		elsif(c = "00110111")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10010010";
			seg3 <= "11000000";
		elsif(c = "00111000")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10010010";
			seg3 <= "11000000";
		elsif(c = "00111001")then	-- 7
			seg1 <= "11111000";
			seg2 <= "10010010";
			seg3 <= "11000000";
		elsif(c = "00111010")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10010010";
			seg3 <= "11000000";
		elsif(c = "00111011")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10010010";
			seg3 <= "11000000";
		elsif(c = "00111100")then	-- 0	60 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "10000010";
			seg3 <= "11000000";
		elsif(c = "00111101")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10000010";
			seg3 <= "11000000";
		elsif(c = "00111110")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10000010";
			seg3 <= "11000000";
		elsif(c = "00111111")then	-- 3 
			seg1 <= "10110000";
			seg2 <= "10000010";
			seg3 <= "11000000";
		elsif(c = "01000000")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10000010";
			seg3 <= "11000000";
		elsif(c = "01000001")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10000010";
			seg3 <= "11000000";
		elsif(c = "01000010")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10000010";
			seg3 <= "11000000";
		elsif(c = "01000011")then	-- 7
			seg1 <= "11111000";
			seg2 <= "10000010";
			seg3 <= "11000000";
		elsif(c = "01000100")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10000010";
			seg3 <= "11000000";
		elsif(c = "01000101")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10000010";
			seg3 <= "11000000";
		elsif(c = "01000110")then	-- 0	70 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "11111000";
			seg3 <= "11000000";
		elsif(c = "01000111")then	-- 1
			seg1 <= "11111001";
			seg2 <= "11111000";
			seg3 <= "11000000";
		elsif(c = "01001000")then	-- 2
			seg1 <= "10100100";
			seg2 <= "11111000";
			seg3 <= "11000000";
		elsif(c = "01001001")then	-- 3
			seg1 <= "10110000";
			seg2 <= "11111000";
			seg3 <= "11000000";
		elsif(c = "01001010")then	-- 4
			seg1 <= "10011001";
			seg2 <= "11111000";
			seg3 <= "11000000";
		elsif(c = "01001011")then	-- 5
			seg1 <= "10010010";
			seg2 <= "11111000";
			seg3 <= "11000000";
		elsif(c = "01001100")then	-- 6
			seg1 <= "10000010";
			seg2 <= "11111000";
			seg3 <= "11000000";
		elsif(c = "01001101")then	-- 7
			seg1 <= "11111000";
			seg2 <= "11111000";
			seg3 <= "11000000";
		elsif(c = "01001110")then	-- 8
			seg1 <= "10000000";
			seg2 <= "11111000";
			seg3 <= "11000000";
		elsif(c = "01001111")then	-- 9
			seg1 <= "10010000";
			seg2 <= "11111000";
			seg3 <= "11000000";
		elsif(c = "01010000")then	-- 0	80 ------------------------------------------- 
			seg1 <= "11000000";	
			seg2 <= "10000000";
			seg3 <= "11000000";
		elsif(c = "01010001")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10000000";
			seg3 <= "11000000";
		elsif(c = "01010010")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10000000";
			seg3 <= "11000000";
		elsif(c = "01010011")then	-- 3	
			seg1 <= "10110000";
			seg2 <= "10000000";
			seg3 <= "11000000";
		elsif(c = "01010100")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10000000";
			seg3 <= "11000000";
		elsif(c = "01010101")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10000000";
			seg3 <= "11000000";
		elsif(c = "01010110")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10000000";
			seg3 <= "11000000";
		elsif(c = "01010111")then	-- 7
			seg1 <= "11111000";
			seg2 <= "10000000";
			seg3 <= "11000000";
		elsif(c = "01011000")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10000000";
			seg3 <= "11000000";
		elsif(c = "01011001")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10000000";
			seg3 <= "11000000";
		elsif(c = "01011010")then	-- 0	90 ------------------------------------------- 
			seg1 <= "11000000";	
			seg2 <= "10010000";
			seg3 <= "11000000";
		elsif(c = "01011011")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10010000";
			seg3 <= "11000000";
		elsif(c = "01011100")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10010000";
			seg3 <= "11000000";
		elsif(c = "01011101")then	-- 3
			seg1 <= "10110000";
			seg2 <= "10010000";
			seg3 <= "11000000";
		elsif(c = "01011110")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10010000";
			seg3 <= "11000000";
		elsif(c = "01011111")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10010000";
			seg3 <= "11000000";
		elsif(c = "01100000")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10010000";
			seg3 <= "11000000";
		elsif(c = "01100001")then	-- 7
			seg1 <= "11111000";
			seg2 <= "10010000";
			seg3 <= "11000000";
		elsif(c = "01100010")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10010000";
			seg3 <= "11000000";
		elsif(c = "01100011")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10010000";
			seg3 <= "11000000";				
		elsif(c = "01100100")then	-- 0	100 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "11000000";
			seg3 <= "11111001";
		elsif(c = "01100101")then	-- 1
			seg1 <= "11111001";
			seg2 <= "11000000";
			seg3 <= "11111001";
		elsif(c = "01100110")then	-- 2
			seg1 <= "10100100";
			seg2 <= "11000000";
			seg3 <= "11111001";
		elsif(c = "01100111")then	-- 3
			seg1 <= "10110000";
			seg2 <= "11000000";
			seg3 <= "11111001";
		elsif(c = "01101000")then	-- 4
			seg1 <= "10011001";
			seg2 <= "11000000";
			seg3 <= "11111001";
		elsif(c = "01101001")then	-- 5
			seg1 <= "10010010";
			seg2 <= "11000000";
			seg3 <= "11111001";
		elsif(c = "01101010")then	-- 6
			seg1 <= "10000010";
			seg2 <= "11000000";
			seg3 <= "11111001";
		elsif(c = "01101011")then	-- 7
			seg1 <= "11111000";
			seg2 <= "11000000";
			seg3 <= "11111001";
		elsif(c = "01101100")then	-- 8
			seg1 <= "10000000";
			seg2 <= "11000000";
			seg3 <= "11111001";
		elsif(c = "01101101")then	-- 9
			seg1 <= "10010000";
			seg2 <= "11000000";
			seg3 <= "11111001";
		elsif(c = "01101110")then	-- 0	110 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "11111001";
			seg3 <= "11111001";
		elsif(c = "01101111")then	-- 1
			seg1 <= "11111001";
			seg2 <= "11111001";
			seg3 <= "11111001";
		elsif(c = "01110000")then	-- 2
			seg1 <= "10100100";
			seg2 <= "11111001";
			seg3 <= "11111001";
		elsif(c = "01110001")then	-- 3
			seg1 <= "10110000";
			seg2 <= "11111001";
			seg3 <= "11111001";
		elsif(c = "01110010")then	-- 4
			seg1 <= "10011001";
			seg2 <= "11111001";
			seg3 <= "11111001";
		elsif(c = "01110011")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10010010";
			seg3 <= "11111001";
		elsif(c = "01110100")then	-- 6
			seg1 <= "10000010";
			seg2 <= "11111001";
			seg3 <= "11111001";
		elsif(c = "01110101")then	-- 7
			seg1 <= "11111000";
			seg2 <= "11111001";
			seg3 <= "11111001";
		elsif(c = "01110110")then	-- 8
			seg1 <= "10000000";
			seg2 <= "11111001";
			seg3 <= "11111001";
		elsif(c = "01110111")then	-- 9
			seg1 <= "10010000";
			seg2 <= "11111001";
			seg3 <= "11111001";
		elsif(c = "01111000")then	-- 0	120 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "10100100";
			seg3 <= "11111001";
		elsif(c = "01111001")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10100100";
			seg3 <= "11111001";
		elsif(c = "01111010")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10100100";
			seg3 <= "11111001";
		elsif(c = "01111011")then	-- 3
			seg1 <= "10110000";
			seg2 <= "10100100";
			seg3 <= "11111001";
		elsif(c = "01111100")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10100100";
			seg3 <= "11111001";
		elsif(c = "01111101")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10100100";
			seg3 <= "11111001";
		elsif(c = "01111110")then	-- 6	
			seg1 <= "10000010";
			seg2 <= "10100100";
			seg3 <= "11111001";
		elsif(c = "01111111")then	-- 7	
			seg1 <= "11111000";
			seg2 <= "10100100";
			seg3 <= "11111001";
		elsif(c = "10000000")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10100100";
			seg3 <= "11111001";
		elsif(c = "10000001")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10100100";
			seg3 <= "11111001";
		elsif(c = "10000010")then	-- 0	130 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "10110000";
			seg3 <= "11111001";
		elsif(c = "10000011")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10110000";
			seg3 <= "11111001";
		elsif(c = "10000100")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10110000";
			seg3 <= "11111001";
		elsif(c = "10000101")then	-- 3
			seg1 <= "10110000";
			seg2 <= "10110000";
			seg3 <= "11111001";
		elsif(c = "10000110")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10110000";
			seg3 <= "11111001";
		elsif(c = "10000111")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10110000";
			seg3 <= "11111001";
		elsif(c = "10001000")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10110000";
			seg3 <= "11111001";
		elsif(c = "10001001")then	-- 7
			seg1 <= "11111000";
			seg2 <= "10110000";
			seg3 <= "11111001";
		elsif(c = "10001010")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10110000";
			seg3 <= "11111001";
		elsif(c = "10001011")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10110000";
			seg3 <= "11111001";
		elsif(c = "10001100")then	-- 0	140 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "10011001";
			seg3 <= "11111001";
		elsif(c = "10001101")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10011001";
			seg3 <= "11111001";
		elsif(c = "10001110")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10011001";
			seg3 <= "11111001";
		elsif(c = "10001111")then	-- 3	
			seg1 <= "10110000";
			seg2 <= "10011001";
			seg3 <= "11111001";
		elsif(c = "10010000")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10011001";
			seg3 <= "11111001";
		elsif(c = "10010001")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10011001";
			seg3 <= "11111001";
		elsif(c = "10010010")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10011001";
			seg3 <= "11111001";
		elsif(c = "10010011")then	-- 7
			seg1 <= "11111000";
			seg2 <= "10011001";
			seg3 <= "11111001";
		elsif(c = "10010100")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10011001";
			seg3 <= "11111001";
		elsif(c = "10010101")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10011001";
			seg3 <= "11111001";				
		elsif(c = "10010110")then	-- 0	150 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "10010010";
			seg3 <= "11111001";
		elsif(c = "10010111")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10010010";
			seg3 <= "11111001";
		elsif(c = "10011000")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10010010";
			seg3 <= "11111001";
		elsif(c = "10011001")then	-- 3
			seg1 <= "10110000";
			seg2 <= "10010010";
			seg3 <= "11111001";
		elsif(c = "10011010")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10010010";
			seg3 <= "11111001";
		elsif(c = "10011011")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10010010";
			seg3 <= "11111001";
		elsif(c = "10011100")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10010010";
			seg3 <= "11111001";
		elsif(c = "10011101")then	-- 7
			seg1 <= "11111000";
			seg2 <= "10010010";
			seg3 <= "11111001";
		elsif(c = "10011110")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10010010";
			seg3 <= "11111001";
		elsif(c = "10011111")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10010010";
			seg3 <= "11111001";
		elsif(c = "10100000")then	-- 0	160 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "10000010";
			seg3 <= "11111001";
		elsif(c = "10100001")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10000010";
			seg3 <= "11111001";
		elsif(c = "10100010")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10000010";
			seg3 <= "11111001";
		elsif(c = "10100011")then	-- 3
			seg1 <= "10110000";
			seg2 <= "10000010";
			seg3 <= "11111001";
		elsif(c = "10100100")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10000010";
			seg3 <= "11111001";
		elsif(c = "10100101")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10000010";
			seg3 <= "11111001";
		elsif(c = "10100110")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10000010";
			seg3 <= "11111001";
		elsif(c = "10100111")then	-- 7
			seg1 <= "11111000";
			seg2 <= "10000010";
			seg3 <= "11111001";
		elsif(c = "10101000")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10000010";
			seg3 <= "11111001";
		elsif(c = "10101001")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10000010";
			seg3 <= "11111001";
		elsif(c = "10101010")then	-- 0	170 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "11111000";
			seg3 <= "11111001";
		elsif(c = "10101011")then	-- 1
			seg1 <= "11111001";
			seg2 <= "11111000";
			seg3 <= "11111001";
		elsif(c = "10101100")then	-- 2
			seg1 <= "10100100";
			seg2 <= "11111000";
			seg3 <= "11111001";
		elsif(c = "10101101")then	-- 3
			seg1 <= "10110000";
			seg2 <= "11111000";
			seg3 <= "11111001";
		elsif(c = "10101110")then	-- 4
			seg1 <= "10011001";
			seg2 <= "11111000";
			seg3 <= "11111001";
		elsif(c = "10101111")then	-- 5	
			seg1 <= "10010010";
			seg2 <= "11111000";
			seg3 <= "11111001";
		elsif(c = "10110000")then	-- 6
			seg1 <= "10000010";
			seg2 <= "11111000";
			seg3 <= "11111001";
		elsif(c = "10110001")then	-- 7
			seg1 <= "11111000";
			seg2 <= "11111000";
			seg3 <= "11111001";
		elsif(c = "10110010")then	-- 8
			seg1 <= "10000000";
			seg2 <= "11111000";
			seg3 <= "11111001";
		elsif(c = "10110011")then	-- 9
			seg1 <= "10010000";
			seg2 <= "11111000";
			seg3 <= "11111001";
		elsif(c = "10110100")then	-- 0	180 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "10000000";
			seg3 <= "11111001";
		elsif(c = "10110101")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10000000";
			seg3 <= "11111001";
		elsif(c = "10110110")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10000000";
			seg3 <= "11111001";
		elsif(c = "10110111")then	-- 3
			seg1 <= "10110000";
			seg2 <= "10000000";
			seg3 <= "11111001";
		elsif(c = "10111000")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10000000";
			seg3 <= "11111001";
		elsif(c = "10111001")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10000000";
			seg3 <= "11111001";
		elsif(c = "10111010")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10000000";
			seg3 <= "11111001";
		elsif(c = "10111011")then	-- 7
			seg1 <= "11111000";
			seg2 <= "10000000";
			seg3 <= "11111001";
		elsif(c = "10111100")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10000000";
			seg3 <= "11111001";
		elsif(c = "10111101")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10000000";
			seg3 <= "11111001";
		elsif(c = "10111110")then	-- 0	190 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "10010000";
			seg3 <= "11111001";
		elsif(c = "10111111")then	-- 1	
			seg1 <= "11111001";
			seg2 <= "10010000";
			seg3 <= "11111001";
		elsif(c = "11000000")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10010000";
			seg3 <= "11111001";
		elsif(c = "11000001")then	-- 3
			seg1 <= "10110000";
			seg2 <= "10010000";
			seg3 <= "11111001";
		elsif(c = "11000010")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10010000";
			seg3 <= "11111001";
		elsif(c = "11000011")then	-- 5
			seg1 <= "10010010";
			seg2 <= "10010000";
			seg3 <= "11111001";
		elsif(c = "11000100")then	-- 6
			seg1 <= "10000010";
			seg2 <= "10010000";
			seg3 <= "11111001";
		elsif(c = "11000101")then	-- 7
			seg1 <= "11111000";
			seg2 <= "10010000";
			seg3 <= "11111001";
		elsif(c = "11000110")then	-- 8
			seg1 <= "10000000";
			seg2 <= "10010000";
			seg3 <= "11111001";
		elsif(c = "11000111")then	-- 9
			seg1 <= "10010000";
			seg2 <= "10010000";
			seg3 <= "11111001";								
		elsif(c = "11001000")then	-- 0	200 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "11000000";
			seg3 <= "10100100";
		elsif(c = "11001001")then	-- 1
			seg1 <= "11111001";
			seg2 <= "11000000";
			seg3 <= "10100100";
		elsif(c = "11001010")then	-- 2
			seg1 <= "10100100";
			seg2 <= "11000000";
			seg3 <= "10100100";
		elsif(c = "11001011")then	-- 3
			seg1 <= "10110000";
			seg2 <= "11000000";
			seg3 <= "10100100";
		elsif(c = "11001100")then	-- 4
			seg1 <= "10011001";
			seg2 <= "11000000";
			seg3 <= "10100100";
		elsif(c = "11001101")then	-- 5
			seg1 <= "10010010";
			seg2 <= "11000000";
			seg3 <= "10100100";
		elsif(c = "11001110")then	-- 6
			seg1 <= "10000010";
			seg2 <= "11000000";
			seg3 <= "10100100";
		elsif(c = "11001111")then	-- 7
			seg1 <= "11111000";
			seg2 <= "11000000";
			seg3 <= "10100100";
		elsif(c = "11010000")then	-- 8
			seg1 <= "10000000";
			seg2 <= "11000000";
			seg3 <= "10100100";
		elsif(c = "11010001")then	-- 9
			seg1 <= "10010000";
			seg2 <= "11000000";
			seg3 <= "10100100";
		elsif(c = "11010010")then	-- 0	210 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "11111001";
			seg3 <= "10100100";
		elsif(c = "11010011")then	-- 1
			seg1 <= "11111001";
			seg2 <= "11111001";
			seg3 <= "10100100";
		elsif(c = "11010100")then	-- 2
			seg1 <= "10100100";
			seg2 <= "11111001";
			seg3 <= "10100100";
		elsif(c = "11010101")then	-- 3
			seg1 <= "10110000";
			seg2 <= "11111001";
			seg3 <= "10100100";
		elsif(c = "11010110")then	-- 4
			seg1 <= "10011001";
			seg2 <= "11111001";
			seg3 <= "10100100";
		elsif(c = "11010111")then	-- 5
			seg1 <= "10010010";
			seg2 <= "11111001";
			seg3 <= "10100100";
		elsif(c = "11011000")then	-- 6
			seg1 <= "10000010";
			seg2 <= "11111001";
			seg3 <= "10100100";
		elsif(c = "11011001")then	-- 7
			seg1 <= "11111000";
			seg2 <= "11111001";
			seg3 <= "10100100";
		elsif(c = "11011010")then	-- 8
			seg1 <= "10000000";
			seg2 <= "11111001";
			seg3 <= "10100100";
		elsif(c = "11011011")then	-- 9
			seg1 <= "10010000";
			seg2 <= "11111001";
			seg3 <= "10100100";			
		elsif(c = "11011100")then	-- 0 220 -------------------------------------------
			seg1 <= "11000000";	
			seg2 <= "10100100";
			seg3 <= "10100100";
		elsif(c = "11011101")then	-- 1
			seg1 <= "11111001";
			seg2 <= "10100100";
			seg3 <= "10100100";
		elsif(c = "11011110")then	-- 2
			seg1 <= "10100100";
			seg2 <= "10100100";
			seg3 <= "10100100";
		elsif(c = "11011111")then	-- 3
			seg1 <= "10110000";
			seg2 <= "10100100";
			seg3 <= "10100100";
		elsif(c = "11100000")then	-- 4
			seg1 <= "10011001";
			seg2 <= "10100100";
			seg3 <= "10100100";					
		elsif(c = "11100001")then	-- 225 -------------------------------------------
			seg1 <= "10010010";
			seg2 <= "10100100";
			seg3 <= "10100100";
			
		end if; -- fin du if
	end process; --fin du process

end behavioral;

------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------